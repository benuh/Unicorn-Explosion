module audio_engine(input CLK100MHZ, input jump, input isdead, output audio);

